/*
You are given a module my_dff with two inputs and one output (that implements a D flip-flop). 
Instantiate three of them, then chain them together to make a shift register of length 3. 
The clk port needs to be connected to all instances.
*/

module top_module ( input clk, input d, output q );
    
  wire wire1,wire2;
    
  my_dff uut1 ( .clk(clk) , .d(d) , .q(wire1));
  my_dff uut2 ( .clk(clk) , .d(wire1) , .q(wire2));
  my_dff uut3 ( .clk(clk) , .d(wire2) , .q(q));
    
endmodule
